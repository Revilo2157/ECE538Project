module large_not(out, A);
        
    input [31:0] A;
    output [31:0] out;

    not or_0(out[0],A[0]);
    not or_1(out[1],A[1]);
    not or_2(out[2],A[2]);
    not or_3(out[3],A[3]);
    not and_4(out[4],A[4]);
    not and_5(out[5],A[5]);
    not and_6(out[6],A[6]);
    not and_7(out[7],A[7]);
    not and_8(out[8],A[8]);
    not and_9(out[9],A[9]);
    not and_10(out[10],A[10]);
    not and_11(out[11],A[11]);
    not and_12(out[12],A[12]);
    not and_13(out[13],A[13]);
    not and_14(out[14],A[14]);
    not and_15(out[15],A[15]);
    not and_16(out[16],A[16]);
    not and_17(out[17],A[17]);
    not and_18(out[18],A[18]);
    not and_19(out[19],A[19]);
    not and_20(out[20],A[20]);
    not and_21(out[21],A[21]);
    not and_22(out[22],A[22]);
    not and_23(out[23],A[23]);
    not and_24(out[24],A[24]);
    not and_25(out[25],A[25]);
    not and_26(out[26],A[26]);
    not and_27(out[27],A[27]);
    not and_28(out[28],A[28]);
    not and_29(out[29],A[29]);
    not and_30(out[30],A[30]);
    not and_31(out[31],A[31]);

endmodule