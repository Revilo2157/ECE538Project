module register_65 (out, in, clk, en, out_en, clr);
   
    input clk, en, clr, out_en;
    input[64:0] in;

    output[64:0] out;

    wire[64:0] dffe_out;

    dffe_ref d0(dffe_out[0],in[0],clk,en,clr);
    dffe_ref d1(dffe_out[1],in[1],clk,en,clr);
    dffe_ref d2(dffe_out[2],in[2],clk,en,clr);
    dffe_ref d3(dffe_out[3],in[3],clk,en,clr);
    dffe_ref d4(dffe_out[4],in[4],clk,en,clr);
    dffe_ref d5(dffe_out[5],in[5],clk,en,clr);
    dffe_ref d6(dffe_out[6],in[6],clk,en,clr);
    dffe_ref d7(dffe_out[7],in[7],clk,en,clr);
    dffe_ref d8(dffe_out[8],in[8],clk,en,clr);
    dffe_ref d9(dffe_out[9],in[9],clk,en,clr);
    dffe_ref d10(dffe_out[10],in[10],clk,en,clr);
    dffe_ref d11(dffe_out[11],in[11],clk,en,clr);
    dffe_ref d12(dffe_out[12],in[12],clk,en,clr);
    dffe_ref d13(dffe_out[13],in[13],clk,en,clr);
    dffe_ref d14(dffe_out[14],in[14],clk,en,clr);
    dffe_ref d15(dffe_out[15],in[15],clk,en,clr);
    dffe_ref d16(dffe_out[16],in[16],clk,en,clr);
    dffe_ref d17(dffe_out[17],in[17],clk,en,clr);
    dffe_ref d18(dffe_out[18],in[18],clk,en,clr);
    dffe_ref d19(dffe_out[19],in[19],clk,en,clr);
    dffe_ref d20(dffe_out[20],in[20],clk,en,clr);
    dffe_ref d21(dffe_out[21],in[21],clk,en,clr);
    dffe_ref d22(dffe_out[22],in[22],clk,en,clr);
    dffe_ref d23(dffe_out[23],in[23],clk,en,clr);
    dffe_ref d24(dffe_out[24],in[24],clk,en,clr);
    dffe_ref d25(dffe_out[25],in[25],clk,en,clr);
    dffe_ref d26(dffe_out[26],in[26],clk,en,clr);
    dffe_ref d27(dffe_out[27],in[27],clk,en,clr);
    dffe_ref d28(dffe_out[28],in[28],clk,en,clr);
    dffe_ref d29(dffe_out[29],in[29],clk,en,clr);
    dffe_ref d30(dffe_out[30],in[30],clk,en,clr);
    dffe_ref d31(dffe_out[31],in[31],clk,en,clr);
    dffe_ref d32(dffe_out[32],in[32],clk,en,clr);
    dffe_ref d33(dffe_out[33],in[33],clk,en,clr);
    dffe_ref d34(dffe_out[34],in[34],clk,en,clr);
    dffe_ref d35(dffe_out[35],in[35],clk,en,clr);
    dffe_ref d36(dffe_out[36],in[36],clk,en,clr);
    dffe_ref d37(dffe_out[37],in[37],clk,en,clr);
    dffe_ref d38(dffe_out[38],in[38],clk,en,clr);
    dffe_ref d39(dffe_out[39],in[39],clk,en,clr);
    dffe_ref d40(dffe_out[40],in[40],clk,en,clr);
    dffe_ref d41(dffe_out[41],in[41],clk,en,clr);
    dffe_ref d42(dffe_out[42],in[42],clk,en,clr);
    dffe_ref d43(dffe_out[43],in[43],clk,en,clr);
    dffe_ref d44(dffe_out[44],in[44],clk,en,clr);
    dffe_ref d45(dffe_out[45],in[45],clk,en,clr);
    dffe_ref d46(dffe_out[46],in[46],clk,en,clr);
    dffe_ref d47(dffe_out[47],in[47],clk,en,clr);
    dffe_ref d48(dffe_out[48],in[48],clk,en,clr);
    dffe_ref d49(dffe_out[49],in[49],clk,en,clr);
    dffe_ref d50(dffe_out[50],in[50],clk,en,clr);
    dffe_ref d51(dffe_out[51],in[51],clk,en,clr);
    dffe_ref d52(dffe_out[52],in[52],clk,en,clr);
    dffe_ref d53(dffe_out[53],in[53],clk,en,clr);
    dffe_ref d54(dffe_out[54],in[54],clk,en,clr);
    dffe_ref d55(dffe_out[55],in[55],clk,en,clr);
    dffe_ref d56(dffe_out[56],in[56],clk,en,clr);
    dffe_ref d57(dffe_out[57],in[57],clk,en,clr);
    dffe_ref d58(dffe_out[58],in[58],clk,en,clr);
    dffe_ref d59(dffe_out[59],in[59],clk,en,clr);
    dffe_ref d60(dffe_out[60],in[60],clk,en,clr);
    dffe_ref d61(dffe_out[61],in[61],clk,en,clr);
    dffe_ref d62(dffe_out[62],in[62],clk,en,clr);
    dffe_ref d63(dffe_out[63],in[63],clk,en,clr);
    dffe_ref d64(dffe_out[64],in[64],clk,en,clr);



    tri_state_buff t0(out[0],dffe_out[0],out_en);
    tri_state_buff t1(out[1],dffe_out[1],out_en);
    tri_state_buff t2(out[2],dffe_out[2],out_en);
    tri_state_buff t3(out[3],dffe_out[3],out_en);
    tri_state_buff t4(out[4],dffe_out[4],out_en);
    tri_state_buff t5(out[5],dffe_out[5],out_en);
    tri_state_buff t6(out[6],dffe_out[6],out_en);
    tri_state_buff t7(out[7],dffe_out[7],out_en);
    tri_state_buff t8(out[8],dffe_out[8],out_en);
    tri_state_buff t9(out[9],dffe_out[9],out_en);
    tri_state_buff t10(out[10],dffe_out[10],out_en);
    tri_state_buff t11(out[11],dffe_out[11],out_en);
    tri_state_buff t12(out[12],dffe_out[12],out_en);
    tri_state_buff t13(out[13],dffe_out[13],out_en);
    tri_state_buff t14(out[14],dffe_out[14],out_en);
    tri_state_buff t15(out[15],dffe_out[15],out_en);
    tri_state_buff t16(out[16],dffe_out[16],out_en);
    tri_state_buff t17(out[17],dffe_out[17],out_en);
    tri_state_buff t18(out[18],dffe_out[18],out_en);
    tri_state_buff t19(out[19],dffe_out[19],out_en);
    tri_state_buff t20(out[20],dffe_out[20],out_en);
    tri_state_buff t21(out[21],dffe_out[21],out_en);
    tri_state_buff t22(out[22],dffe_out[22],out_en);
    tri_state_buff t23(out[23],dffe_out[23],out_en);
    tri_state_buff t24(out[24],dffe_out[24],out_en);
    tri_state_buff t25(out[25],dffe_out[25],out_en);
    tri_state_buff t26(out[26],dffe_out[26],out_en);
    tri_state_buff t27(out[27],dffe_out[27],out_en);
    tri_state_buff t28(out[28],dffe_out[28],out_en);
    tri_state_buff t29(out[29],dffe_out[29],out_en);
    tri_state_buff t30(out[30],dffe_out[30],out_en);
    tri_state_buff t31(out[31],dffe_out[31],out_en);
    tri_state_buff t32(out[32],dffe_out[32],out_en);
    tri_state_buff t33(out[33],dffe_out[33],out_en);
    tri_state_buff t34(out[34],dffe_out[34],out_en);
    tri_state_buff t35(out[35],dffe_out[35],out_en);
    tri_state_buff t36(out[36],dffe_out[36],out_en);
    tri_state_buff t37(out[37],dffe_out[37],out_en);
    tri_state_buff t38(out[38],dffe_out[38],out_en);
    tri_state_buff t39(out[39],dffe_out[39],out_en);
    tri_state_buff t40(out[40],dffe_out[40],out_en);
    tri_state_buff t41(out[41],dffe_out[41],out_en);
    tri_state_buff t42(out[42],dffe_out[42],out_en);
    tri_state_buff t43(out[43],dffe_out[43],out_en);
    tri_state_buff t44(out[44],dffe_out[44],out_en);
    tri_state_buff t45(out[45],dffe_out[45],out_en);
    tri_state_buff t46(out[46],dffe_out[46],out_en);
    tri_state_buff t47(out[47],dffe_out[47],out_en);
    tri_state_buff t48(out[48],dffe_out[48],out_en);
    tri_state_buff t49(out[49],dffe_out[49],out_en);
    tri_state_buff t50(out[50],dffe_out[50],out_en);
    tri_state_buff t51(out[51],dffe_out[51],out_en);
    tri_state_buff t52(out[52],dffe_out[52],out_en);
    tri_state_buff t53(out[53],dffe_out[53],out_en);
    tri_state_buff t54(out[54],dffe_out[54],out_en);
    tri_state_buff t55(out[55],dffe_out[55],out_en);
    tri_state_buff t56(out[56],dffe_out[56],out_en);
    tri_state_buff t57(out[57],dffe_out[57],out_en);
    tri_state_buff t58(out[58],dffe_out[58],out_en);
    tri_state_buff t59(out[59],dffe_out[59],out_en);
    tri_state_buff t60(out[60],dffe_out[60],out_en);
    tri_state_buff t61(out[61],dffe_out[61],out_en);
    tri_state_buff t62(out[62],dffe_out[62],out_en);
    tri_state_buff t63(out[63],dffe_out[63],out_en);
    tri_state_buff t64(out[64],dffe_out[64],out_en);


    

endmodule